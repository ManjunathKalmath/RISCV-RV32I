module ALU_Control(ALU_OP,funct_code,ALU_Ctl);
input [1:0] ALU_OP;
input [5:0] funct_code;
Output reg [3:0] ALU_Ctl;

always begin
case (funct_code)
32 : 
end
endmodule
