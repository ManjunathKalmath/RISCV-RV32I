module RV32IM_Controlpath(clock);
  input clock;
endmodule
