module RV32IM_Controlpath(clock);
  input clock;
  //Instantiate ALU_Control here
endmodule
